../lfsr_prnd/lfsr_prnd.vhd