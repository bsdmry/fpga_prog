../spi_slave_drv/spi_slave_drv.vhd