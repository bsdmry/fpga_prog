../uart/uart.vhd