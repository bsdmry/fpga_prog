../mseg_ctl/mseg_ctl.vhd