../ws1228_driver/ws1228_driver.vhd