../dram_ctl/dram_ctl.vhd