../max98257_driver/max98257_driver.vhd